.include 'solar_cell.txt'
 
x1 1 2 solar_cell
vsolar 3 1 dc 0
r1 2 3 100

.dc r1 0.001 10k 0.1
.control

run
let power = {i(vsolar)*(v(1) - v(2))}
let id = i(vsolar)
let vd = {v(1) - v(2)}
plot id vs vd power vs vd  
.endc
.end
