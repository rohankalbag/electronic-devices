*IV Characteristics
*Rohan Rajesh Kalbag 20D170033
.include yellow_5mm.txt
.include red_5mm.txt
.include green_5mm.txt
.include blue_5mm.txt
.include white_5mm.txt
.include Diode_1N914.txt

vs 1 0 dc 0

vyellow 21 31 dc 0
da 1 21 YELLOW
ra 31 0 100

vred 22 32 dc 0
db 1 22 RED
rb 32 0 100

vgreen 23 33 dc 0
dc 1 23 GREEN
rc 33 0 100

vblue 24 34 dc 0
dd 1 24 BLUE
rd 34 0 100

vwhite 25 35 dc 0
de 1 25 WHITE
re 35 0 100

v1n914 26 36 dc 0
df 1 26 1N914
rf 36 0 100

.dc vs 0.001 5 0.01
.control

run
plot i(vyellow) vs v(1) - v(21) i(vred) vs v(1) - v(22) i(vgreen) vs v(1) - v(23) i(vblue) vs v(1) - v(24) i(vwhite) vs v(1) - v(25) i(v1n914) vs v(1) - v(26)
plot ln(i(vyellow)) vs v(1) - v(21) ln(i(vred)) vs v(1) - v(22) ln(i(vgreen)) vs v(1) - v(23) ln(i(vblue)) vs v(1) - v(24) ln(i(vwhite)) vs v(1) - v(25) ln(i(v1n914)) vs v(1) - v(26)
.endc
.end