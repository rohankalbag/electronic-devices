Forward Voltage and Current for varying Temperature 

.include 'photo_diode.txt'

v1 0 1 -1.5 dc 
x1 1 2 photo_diode IL_val=1e-3
vdiode 2 3 dc 0
r1 3 0 100

.op
.option set temp = 75
.control

run
print i(vdiode)
print v(1) - v(2)
.endc
.end
