Dark IV Characteristics 1(a)

.include 'photo_diode.txt'

v1 0 1 dc 
x1 1 2 photo_diode IL_val=0e-3
vdiode 2 3 dc 0
r1 3 0 100

.dc v1 -2 2 0.01
.control

run
let id = i(vdiode)
let vd = {v(1) - v(2)}
plot id vs vd
.endc
.end
